module top();

endmodule top();