module registerfile();

endmodule registerfile();