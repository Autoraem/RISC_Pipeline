module regfile();

endmodule regfile();